`include alu_controll.vh
`include Opcode.vh

module alu_controller(
	input [31:0] instruction,
	output [3:0] alu_controll
	);

wire [6:0] opcode;
assign opcode = instruction[6:0];

wire [2:0] funct3;
assign funct3 = instruction[14:12];

wire [6:0] funct7;
assign funct7 = instruction[31:25];


always @(*) begin
	case(opcode)
		OPC_ARI_RTYPE: begin
							case(funct3)
								3'b000: begin
									case(funct7)
										7'b0000000: alu_controll = ADD;
										7'b0100000: alu_controll = SUB;
										default: begin
											alu_controll = NOP;
											$display("Undefined instruction in alu_controller");
										end
									endcase
								end
								3'b001: alu_controll = SLL;
								3'b010: alu_controll = LT;
								3'b011: alu_controll = LTU;
								3'b100: alu_controll = XOR;
								3'b101: begin
									case(funct7)
										7'b0000000: alu_controll = SRL;
										7'b0100000: alu_controll = SRA;
										default: begin
											alu_controll = NOP;
											$display("Undefined instruction in alu_controller");
										end
									endcase
								end
								3'b110: alu_controll = OR;
								3'b111: alu_controll = AND;
							endcase
					   end
		OPC_ARI_ITYPE: begin
							case(funct3)
								3'b000: alu_controll = ADD;
								3'b001: alu_controll = SLL;
								3'b010: alu_controll = LT;
								3'b011: alu_controll = LTU;
								3'b100: alu_controll = XOR;
								3'b101: begin
									case(funct7)
										7'b0000000: alu_controll = SRL;
										7'b0100000: alu_controll = SRA;
										default: begin
											alu_controll = NOP;
											$display("Undefined instruction in alu_controller");
										end
									endcase
								end
								3'b110: alu_controll = OR;
								3'b111: alu_controll = AND;
							endcase
					   end
		OPC_LOAD:  alu_controll = ADD;
		OPC_STORE: alu_controll = ADD;
		OPC_JALR:  alu_controll = ADD;
		OPC_JAL: begin
					alu_controll = NOP;
					$display("JAL in alu_controller");
				 end
		OPC_BRANCH: alu_controller = SUB;
		OPC_AUIPC:  alu_controller = ADD;
		OPC_LUI:	alu_controller = NOP; // No ALU operation needed
	endcase
end


endmodule