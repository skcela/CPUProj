`include "mux_selects.vh"
`include "Opcode.vh"
/**
 * Top-level module for the RISCV processor.
 * Contains instantiations of datapath and control unit.
 */
module Riscv151 #(
    parameter CPU_CLOCK_FREQ = 50_000_000
)(
    input clk,
    input rst,

    output io_fifo_rd_en,
    input [7:0] io_fifo_dout,
    input io_fifo_empty,

    input [7:0] gpio_switches,

    output [12:0] leds_dout,

    output tone_generator_enable,
    output [23:0] tone_generator_switch_period,

    input ac_fifo_full,
    output ac_fifo_wr_en,
    output [19:0] ac_fifo_din,
    output [3:0] ac_volume,

    input mic_fifo_empty,
    output mic_fifo_read_en,
    input [31:0] mic_fifo_dout,

    // Ports for i2c
    input [15:0] i2c_rdata,

    output [15:0] i2c_wdata_unreg,
    output [15:0] i2c_slave_addr_unreg,
    output [15:0] i2c_reg_addr_unreg,

    input i2c_ctrl_ready,
    output i2c_ctrl_valid,

    output i2c_rdata_ready,
    input i2c_rdata_valid,

    output arb_we,
    output arb_din,
    output [19:0] arb_addr,

    // Ports for UART that go off-chip to UART level shifter
    input FPGA_SERIAL_RX,
    output FPGA_SERIAL_TX
);


    // ------------------------- Connections for PC / Instruction -------------------------
    // Pipeline registers for pc in different stages
    reg [31:0] pc;
    wire [31:0] pc_plus_4;
    reg [31:0] next_pc;
    assign pc_plus_4 = pc + 4;
    reg [31:0] pc_2;
    reg [31:0] pc_3;
    reg [31:0] pc_plus_4_2;
    reg [31:0] pc_plus_4_3;
    always @(posedge clk) begin
        pc_2 <= pc;
        pc_3 <= pc_2;
        pc_plus_4_2 <= pc_plus_4;
        pc_plus_4_3 <= pc_plus_4_2;
    end
    // Reset of PC
    always @(posedge clk) begin
        if (rst) begin
            // reset
            pc <= 32'h3FFFFFFC;
        end
        else begin
            pc <= next_pc;
        end
    end

    // Instruction in first stage
    wire [31:0] bios_mem_instruction_out;
    wire [31:0] imem_instruction_out;
    wire [31:0] instruction_1;
    assign instruction_1 =  (pc == 32'h3FFFFFFC) ? 32'b0  :
                                          pc[30] ? bios_mem_instruction_out 
                                                 : imem_instruction_out;
    // Instruction in second and third stage, generated by control unit
    wire [31:0] instruction_2;
    wire [31:0] instruction_3;
    wire [6:0] opcode_2;
    assign opcode_2 = instruction_2[6:0];
    wire [6:0] opcode_3;
    assign opcode_3 = instruction_3[6:0];

    // Mux for next pc
    // PC Mux select signal, generated by control unit
    wire [`PC_MUX_SEL_WIDTH-1:0] pc_mux_sel;
    // branch address and alu output as calculated in stage 2
    wire [31:0] branch_address;
    wire [31:0] alu_out;
    always @(*) begin
        case(pc_mux_sel)
            `PC_MUX_BRANCH: next_pc = branch_address;
            `PC_MUX_J:      next_pc = alu_out;
            default:        next_pc = pc_plus_4;
        endcase
    end


    // ------------------------- Connections for CONTROLLUNIT -------------------------   
    wire [`WB_MUX_SEL_WIDTH-1:0] wb_mux_sel;
    wire [`ALU_IN_MUX_SEL_WIDTH-1:0] alu_in_mux_1_sel;
    wire [`ALU_IN_MUX_SEL_WIDTH-1:0] alu_in_mux_2_sel;
    wire branch_condition;
    wire store_wb_hazard;
    wire wb_reg_hazard_rs1;
    wire wb_reg_hazard_rs2;
    // connection from controll unit to mem controller for store hazard
    wire store_alu_hazard;


    // ------------------------- Connections for DATAPATH -------------------------
    // Connections for alu input muxes to alu
    wire [31:0] alu_in_1;
    wire [31:0] alu_in_2;

    // register for alu_out in third pipeline stage
    reg [31:0] alu_out_3;
    always @(posedge clk) begin
        alu_out_3 <= alu_out;
    end

    // connections for reg file
    wire rf_write_enable;
    wire [31:0] rf_write_data;
    wire [31:0] rd1;
    wire [31:0] rd2;
    // pipeline registers for reg file output
    reg [31:0] rd1_2;
    reg [31:0] rd2_2;
    reg [31:0] mem_data_in;
    // Registers for first pipeline stage
    always @(posedge clk ) begin
        rd1_2 <= wb_reg_hazard_rs1 ? rf_write_data : rd1;
        rd2_2 <= wb_reg_hazard_rs2 ? rf_write_data : rd2;
        mem_data_in <= store_wb_hazard ? rf_write_data : rd2;
    end


    // ------------------------- Connections for MEMORIES -------------------------
    wire [3:0] write_enable_mask; // says which byte should be written
    // enable signal for all memories
    wire [3:0] imem_write_enable;
    wire [3:0] dmem_write_enable; 
    wire cycle_counter_write_enable;
    wire uart_write_enable;
    wire led_write_enable;
    // data connections for read and write controller and memories
    wire [31:0] mem_controller_data_out;
    wire [31:0] dmem_data_out;
    wire [31:0] bios_mem_data_out;
    wire [31:0] cycle_counter_dout;
    wire [31:0] mem_dout;
    wire [7:0] uart_dout;
    wire uart_din_ready;
    wire uart_dout_valid;
    wire [31:0] uart_data_0;
    wire [31:0] uart_data_4;
    assign uart_data_0 = {30'b0, uart_dout_valid, uart_din_ready};
    assign uart_data_4 = {24'b0, uart_dout};
    // Ready - Valid interface for UART
    wire uart_dout_ready;
    assign uart_dout_ready = (((alu_out_3 == 32'h80000000) | (alu_out_3 == 32'h80000004))
                              & (opcode_3 == `OPC_LOAD));

    // Read enable for fifo, set in stage 2 becaus it's a synchronous read
    assign io_fifo_rd_en = ((alu_out == 32'h80000024)
                              & (opcode_2 == `OPC_LOAD));


    // Ready - Valid interface for I2C controller
    assign i2c_rdata_ready = ((alu_out_3 == 32'h80000104)
                              & (opcode_3 == `OPC_LOAD));


    // write to tone generator
    reg tone_generator_enable_reg;
    reg [23:0] tone_generator_switch_period_reg;
    assign tone_generator_enable = tone_generator_enable_reg;
    assign tone_generator_switch_period = tone_generator_switch_period_reg;
    always @(posedge clk) begin
        if (rst) begin
            // reset
            tone_generator_enable_reg <= 0;
        end
        else if ((alu_out == 32'h80000034) & (opcode_2 == `OPC_STORE)) begin
            tone_generator_enable_reg <= mem_controller_data_out[0];
        end
    end

    always @(posedge clk) begin
        if (rst) begin
            // reset
            tone_generator_switch_period_reg <= 0;
        end
        else if ((alu_out == 32'h80000038) & (opcode_2 == `OPC_STORE)) begin
            tone_generator_switch_period_reg <= mem_controller_data_out[23:0];
        end
    end

    // write to ac97 controller
    reg [19:0] ac_fifo_din_reg;
    reg [3:0] ac_volume_reg;
    reg ac_fifo_wr_en_reg;
    assign ac_fifo_din = ac_fifo_din_reg;
    assign ac_volume = ac_volume_reg;
    assign ac_fifo_wr_en = ac_fifo_wr_en_reg;
    always @(posedge clk) begin
        if (rst) begin
            // reset
            ac_fifo_din_reg <= 0;
            ac_fifo_wr_en_reg <= 0;
        end
        else if ((alu_out == 32'h80000044) & (opcode_2 == `OPC_STORE)) begin
            ac_fifo_din_reg <= mem_controller_data_out[19:0];
            ac_fifo_wr_en_reg <= 1;
        end else begin
            ac_fifo_wr_en_reg <= 0;
            ac_fifo_din_reg <= 0;
        end
    end

    always @(posedge clk) begin
        if (rst) begin
            // reset
            ac_volume_reg <= 0;
        end
        else if ((alu_out == 32'h80000048) & (opcode_2 == `OPC_STORE)) begin
            ac_volume_reg <= mem_controller_data_out[3:0];
        end
    end

    assign mic_fifo_read_en = ((alu_out == 32'h80000054) & (opcode_2 == `OPC_LOAD));

    // write the LEDs
    reg [12:0] leds_reg;
    assign leds_dout = leds_reg;
    always @(posedge clk) begin
        if (rst) begin
            // reset
            leds_reg <= 0;
        end
        else if (led_write_enable) begin
            leds_reg <= mem_controller_data_out[13:0];
        end
    end


    // Write to i2c controller
    reg [15:0] i2c_reg_addr, i2c_wdata, i2c_slave_addr;
    assign i2c_slave_addr_unreg = i2c_slave_addr;
    assign i2c_wdata_unreg = i2c_wdata;
    assign i2c_reg_addr_unreg = i2c_reg_addr;
    reg i2c_ctrl_valid_reg;
    assign i2c_ctrl_valid = i2c_ctrl_valid_reg;

    always @(posedge clk) begin
        if(rst) begin
            i2c_reg_addr <= 0;
            i2c_wdata <= 0;
            i2c_slave_addr <= 0;
            i2c_ctrl_valid_reg <= 0;
        end else if (opcode_2 == `OPC_STORE) begin
            if (alu_out == 32'h80000108) begin
                i2c_reg_addr <= mem_controller_data_out[15:0];
            end

            if (alu_out == 32'h8000010C) begin
                i2c_wdata <= mem_controller_data_out[15:0];                
            end
            
            if (alu_out == 32'h80000110) begin
                i2c_slave_addr <= mem_controller_data_out[15:0];                
            end

            if (alu_out == 32'h80000114) begin
                i2c_ctrl_valid_reg <= 1;
            end
        end

        if (i2c_ctrl_valid_reg) begin
                i2c_ctrl_valid_reg <= 0;
        end
    end

    // write to frame buffer
    wire frame_buffer_wen;
    reg [19:0] arb_addr_reg;
    assign arb_addr = arb_addr_reg;
    reg arb_din_reg, arb_we_reg;
    assign arb_din = arb_din_reg;
    assign arb_we = arb_we_reg;
    always @(posedge clk) begin
        if (rst) begin
            // reset
            arb_we_reg <= 0;
            arb_addr_reg <= 0;
            arb_din_reg <= 0;
        end
        else if (frame_buffer_wen) begin
            arb_addr_reg <= alu_out[19:0];
            arb_din_reg <= mem_controller_data_out[0];
            arb_we_reg <= 1;
        end else begin
            arb_we_reg <= 0;
            arb_din_reg <= 0;
            arb_addr_reg <= 0;
        end
    end

    // ------------------------------ MEMORIES - I/O ------------------------------
    mem_write_controller mem_write_controller(
        .instruction(instruction_2),
        .address(alu_out),
        .data_in(store_alu_hazard ? rf_write_data :  mem_data_in),
        .data_out(mem_controller_data_out),
        .write_enable_mask(write_enable_mask),
        .dmem_write_enable(dmem_write_enable),
        .imem_write_enable(imem_write_enable),
        .led_write_enable(led_write_enable),
        .cycle_counter_write_enable(cycle_counter_write_enable),
        .uart_write_enable(uart_write_enable),
        .frame_buffer_wen(frame_buffer_wen)
    );

    dmem_blk_ram dmem (
        .clka(clk),
        .ena(1'b1),
        .wea(dmem_write_enable & write_enable_mask),
        .addra(alu_out[15:2]),
        .dina(mem_controller_data_out),
        .douta(dmem_data_out)
    );

    bios_mem bios_mem(
        .clka(clk),
        .clkb(clk),
        .ena(1'b1),
        .enb(1'b1),
        .addra(next_pc[15:2]),
        .douta(bios_mem_instruction_out),
        .addrb(alu_out[15:2]),
        .doutb(bios_mem_data_out)
    );

    imem_blk_ram imem( 
        .clka(clk),
        .clkb(clk),
        .ena(1'b1),
        .wea(imem_write_enable & write_enable_mask),
        .addra(alu_out[15:2]),
        .dina(mem_controller_data_out),
        .addrb(next_pc[15:2]),
        .doutb(imem_instruction_out)
    );

    cycle_counter cycle_counter(
        .clk(clk),
        .rst(rst),
        .instruction_3(instruction_3),
        .address(alu_out),
        .write_enable(cycle_counter_write_enable),
        .d_in(mem_controller_data_out),
        .d_out(cycle_counter_dout)
    );

    mem_read_controller mem_read_controller(
        .instruction(instruction_3),
        .mem_addr(alu_out_3),
        .dmem_data_in(dmem_data_out),
        .bios_data_in(bios_mem_data_out),
        .uart_data_0_in(uart_data_0),
        .uart_data_4_in(uart_data_4),
        .io_fifo_empty(io_fifo_empty),
        .io_fifo_dout(io_fifo_dout),
        .gpio_switches(gpio_switches),
        .cycle_counter_data_in(cycle_counter_dout),
        .ac_fifo_full(ac_fifo_full),
        .mic_fifo_empty(mic_fifo_empty),
        .mic_fifo_dout(mic_fifo_dout),

        .i2c_rdata_valid(i2c_rdata_valid),
        .i2c_ctrl_ready(i2c_ctrl_ready),
        .i2c_rdata(i2c_rdata),

        .data_out(mem_dout)
    );

    // On-chip UART
    uart #(
        .CLOCK_FREQ(CPU_CLOCK_FREQ)
    ) on_chip_uart (
        .clk(clk),
        .reset(rst),
        .data_in(mem_controller_data_out[7:0]),
        .data_in_valid(uart_write_enable),
        .data_out_ready(uart_dout_ready),
        .serial_in(FPGA_SERIAL_RX),

        .data_in_ready(uart_din_ready),
        .data_out(uart_dout),
        .data_out_valid(uart_dout_valid),
        .serial_out(FPGA_SERIAL_TX)
    );


    // ------------------------------ CONTROLL UNIT ------------------------------

    control_unit control_unit(
        .clk(clk),
        .rst(rst),
        .instruction_1(instruction_1),
        .instruction_2_o(instruction_2),
        .instruction_3_o(instruction_3),
        .branch_condition(branch_condition),
        .wb_reg_hazard_rs1(wb_reg_hazard_rs1),
        .wb_reg_hazard_rs2(wb_reg_hazard_rs2),
        .store_alu_hazard(store_alu_hazard),
        .store_wb_hazard(store_wb_hazard),
        .alu_in_mux_1_sel(alu_in_mux_1_sel),
        .alu_in_mux_2_sel(alu_in_mux_2_sel),
        .wb_mux_sel(wb_mux_sel),
        .pc_mux_sel(pc_mux_sel)
    );


    branch_checker branch_checker(
        .instruction_2(instruction_2),
        .alu_output(alu_out),
        .branch_condition(branch_condition)
    );

    // ------------------------------ DATAPATH ------------------------------
    
    reg_file rf(
        .clk(clk),
        .rst(rst),
        .we(rf_write_enable),
        .ra1(instruction_1[19:15]), 
        .ra2(instruction_1[24:20]), 
        .wa(instruction_3[11:7]),
        .wd(rf_write_data),
        .rd1(rd1), 
        .rd2(rd2)
    );

    alu_in_muxes alu_in_muxes(
        .instruction(instruction_2),
        .mux_1_sel(alu_in_mux_1_sel),
        .mux_2_sel(alu_in_mux_2_sel),
        .rd1(rd1_2),
        .rd2(rd2_2),
        .pc(pc_2),
        .fw_writeback(rf_write_data),
        
        .alu_in_1(alu_in_1), 
        .alu_in_2(alu_in_2)
    );

    stage2 stage2(
        .instruction_in(instruction_2),

        .alu_in_1(alu_in_1),
        .alu_in_2(alu_in_2),
        .alu_out(alu_out),

        // pc for calculation of branch address
        .pc(pc_2),
        .branch_address(branch_address)
    );


    writeback_mux writeback_mux(
        .instruction(instruction_3),
        .mux_sel(wb_mux_sel),
        .pc_plus_4(pc_plus_4_3),
        .mem_dout(mem_dout),
        .alu_out(alu_out_3),
        .writeback_data(rf_write_data),
        .writeback_enable(rf_write_enable)
    );





endmodule
